Decimal Hexadecimal Octal Symbol\Char
000 00 000 NUL
001 01 001 SOH
002 02 002 STX
003 03 003 ETX
004 04 004 EOT
005 05 005 ENQ
006 06 006 ACK
007 07 007 BEL
008 08 010 BS
009 09 011 TAB
010 0A 012 NL
011 0B 013 VT
012 0C 014 NP
013 0D 015 CR
014 0E 016 SO
015 0F 017 SI
016 10 020 DLE
017 11 021 DC1
018 12 022 DC2
019 13 023 DC3
020 14 024 DC4
021 15 025 NAK
022 16 026 SYN
023 17 027 ETB
024 18 030 CAN
025 19 031 EM
026 1A 032 SUB
027 1B 033 ESC
028 1C 034 FS
029 1D 035 GS
030 1E 036 RS
031 1F 037 US
032 20 040 SP
033 21 041 !
034 22 042 "
035 23 043 #
036 24 044 $
037 25 045 %
038 26 046 &
039 27 047 '
040 28 050 (
041 29 051 )
042 2A 052 *
043 2B 053 +
044 2C 054 ,
045 2D 055 -
046 2E 056 .
047 2F 057 /
048 30 060 0
049 31 061 1
050 32 062 2
051 33 063 3
052 34 064 4
053 35 065 5
054 36 066 6
055 37 067 7
056 38 070 8
057 39 071 9
058 3A 072 :
059 3B 073 ;
060 3C 074 <
061 3D 075 =
062 3E 076 >
063 3F 077 ?
064 40 100 @
065 41 101 A
066 42 102 B
067 43 103 C
068 44 104 D
069 45 105 E
070 46 106 F
071 47 107 G
072 48 110 H
073 49 111 I
074 4A 112 J
075 4B 113 K
076 4C 114 L
077 4D 115 M
078 4E 116 N
079 4F 117 O
080 50 120 P
081 51 121 Q
082 52 122 R
083 53 123 S
084 54 124 T
085 55 125 U
086 56 126 V
087 57 127 W
088 58 130 X
089 59 131 Y
090 5A 132 Z
091 5B 133 [
092 5C 134 \
093 5D 135 ]
094 5E 136 ^
095 5F 137 _
096 60 140 `
097 61 141 a
098 62 142 b
099 63 143 c
100 64 144 d
101 65 145 e
102 66 146 f
103 67 147 g
104 68 150 h
105 69 151 i
106 6A 152 j
107 6B 153 k
108 6C 154 l
109 6D 155 m
110 6E 156 n
111 6F 157 o
112 70 160 p
113 71 161 q
114 72 162 r
115 73 163 s
116 74 164 t
117 75 165 u
118 76 166 v
119 77 167 w
120 78 170 x
121 79 171 y
122 7A 172 z
123 7B 173 {
124 7C 174 |
125 7D 175 }
126 7E 176 ~
127 7F 177 DEL
